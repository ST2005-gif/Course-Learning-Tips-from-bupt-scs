module v14(
    input [3:0] a, 
    output reg [7:0] y  
);

always @(*) begin
    case (a)
        4'b0000: y = 7'b1111110;//0
        4'b0001: y = 7'b0110000;//1
        4'b0010: y = 7'b1101101;//2
        4'b0011: y = 7'b1111001;//3
        4'b0100: y = 7'b0110011;//4
        4'b0101: y = 7'b1011011;//5
        4'b0110: y = 7'b0011111;//6
        4'b0111: y = 7'b1110000;//7
        4'b1000: y = 7'b1111111;//8
        4'b0111: y = 7'b1110011;//9
        default: y = 7'b0000000;//other
    endcase
end

endmodule